`ifndef _parameters_vh_
`define _parameters_vh_
parameter       maxVert = 524;
parameter       maxHorz = 799;
parameter       syncVert = 2;
parameter       syncHorz = 96;
parameter       activeHorzmax = 784;
parameter       activeHorzmin = 143;
parameter       activeVertmax = 515;
parameter       activeVertmin = 35;
`endif